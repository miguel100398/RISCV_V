//File: riscv_v_alu_scbd.sv
//Author: Miguel Bucio
//Date: 11/06/23
//Description: RISC-V Vector ALU Scoreboard

`ifndef __RISCV_V_ALU_SCBD_SV__
`define __RISCV_V_ALU_SCBD_SV__ 

class riscv_v_alu_scbd extends riscv_v_base_scbd#(
                                                 .seq_item_in_t(riscv_v_alu_in_seq_item),
                                                 .seq_item_out_t(riscv_v_alu_out_seq_item) );
    `uvm_component_utils(riscv_v_alu_scbd)

    riscv_v_logic_alu_in_seq_item       logic_in_txn;
    riscv_v_arithmetic_alu_in_seq_item  arithmetic_in_txn;
    riscv_v_mask_alu_in_seq_item        mask_in_txn;
    riscv_v_permutation_alu_in_seq_item permutation_in_txn;

    //Expected results
    riscv_v_wb_data_t  logic_exp_result;
    riscv_v_wb_data_t  arithmetic_exp_result;
    riscv_v_mask_t     mask_exp_result;
    riscv_v_wb_data_t  permutation_exp_vec_result;
    riscv_data_t       permutation_exp_int_result;
    riscv_v_zf_t       zf_exp;
    riscv_v_of_t       of_exp;
    riscv_v_cf_t       cf_exp;

    function new(string name = "riscv_v_alu_scbd", uvm_component parent = null);
        super.new(name, parent);
    endfunction: new

    virtual function void calc_in();
        //Cast transaction
        calc_valid();
        if ($cast(logic_in_txn, txn_in)) begin
            calc_logic();
        end else if ($cast(arithmetic_in_txn, txn_in))begin
            calc_arithmetic();
        end else if ($cast(mask_in_txn, txn_in)) begin
            calc_mask();
        end else if ($cast(permutation_in_txn, txn_in)) begin 
            calc_permutation();
        end else begin
            `uvm_fatal(get_name(), "Can't cast alu_seq_in to valid specific_alu_seq_in")
        end
    endfunction: calc_in 

    virtual function void calc_out();
        case(txn_out.ALU) 
            LOGIC_ALU: compare_logic();
            ARITHMETIC_ALU: compare_arithmetic();
            MASK_ALU: compare_mask();
            PERMUTATION_ALU: compare_permutation();
            default:   `uvm_fatal(get_name(), "Invalid ALU found in txn_out")
        endcase
    endfunction: calc_out

    virtual function void calc_logic();
        case(logic_in_txn.opcode)
            BW_AND:         calc_bw_and();
            BW_AND_REDUCT:  calc_bw_and_reduct();
            BW_OR:          calc_bw_or();
            BW_OR_REDUCT:   calc_bw_or_reduct();
            BW_XOR:         calc_bw_xor();
            BW_XOR_REDUCT:  calc_bw_xor_reduct();
            SLL:            calc_sll();
            SRL:            calc_srl();
            SRA:            calc_sra();
            default:        `uvm_fatal(get_name(), "Invalid Logic ALU op")
        endcase
    endfunction: calc_logic

    virtual function void calc_arithmetic();
        case(arithmetic_in_txn.opcode)
            ADDC:           calc_addc();
            ADD:            calc_add();
            ADD_REDUCT:     calc_add_reduct();
            SUBB:           calc_subb();
            SUB:            calc_sub();
            SUB_REDUCT:     calc_sub_reduct();
            SIGN_EXT:       calc_sign_ext();
            ZERO_EXT:       calc_zero_ext();
            MINS:           calc_mins();
            MINS_REDUCT:    calc_mins_reduct();
            MINU:           calc_minu();
            MINU_REDUCT:    calc_minu_reduct();
            MAXS:           calc_maxs();
            MAXS_REDUCT:    calc_maxs_reduct();
            MAXU:           calc_maxu();
            MAXU_REDUCT:    calc_maxu_reduct();
            MULLU:          calc_mullu();
            MULLS:          calc_mulls();
            MULHU:          calc_mulhu();
            MULHS:          calc_mulhs();
            SEQ:            calc_seq();
            SNE:            calc_sne();
            SLE:            calc_sle();
            SLEU:           calc_sleu();
            SLT:            calc_slt();
            SLTU:           calc_sltu();
            SGT:            calc_sgt();
            SGTU:           calc_sgtu();
            default:        `uvm_fatal(get_name(), "Invalid arithmetic ALU op")
        endcase
    endfunction: calc_arithmetic

    virtual function void calc_mask();
        case(mask_in_txn.opcode)
            MAND:   calc_mand();
            MNAND:  calc_mnand();
            MANDN:  calc_mandn();
            MOR:    calc_mor();
            MNOR:   calc_mnor();
            MORN:   calc_morn();
            MXOR:   calc_mxor();
            MXNOR:  calc_mxnor();
            default: `uvm_fatal(get_name(), "Invalid mask ALU op")
        endcase
    endfunction: calc_mask

    virtual function void calc_permutation();
        case(permutation_in_txn.opcode)
            I2V: calc_i2v();
            V2I: calc_v2i();
            default: `uvm_fatal(get_name(), "Invalid permutation ALU op")
        endcase
    endfunction: calc_permutation

    virtual function void compare_logic();
        bit comp = 1;
        comp &= logic_exp_result.valid == txn_out.result.valid;
        for (int i=0; i<RISCV_V_NUM_BYTES_DATA; i++) begin
            if (logic_exp_result.valid[i]) begin
                comp &= logic_exp_result.data.Byte[i] == txn_out.result.data.Byte[i];
            end
        end
        if (comp) begin
            pass();
        end else begin
            `uvm_error(get_name(), $sformatf("Compare mismatch, actual.valid: 0x%0h, actual.data 0x%0h, exp.valid: 0x%0h, exp.data: 0x%0h", txn_out.result.valid, txn_out.result.data, logic_exp_result.valid, logic_exp_result.data))
            fail();
        end
    endfunction: compare_logic

    virtual function void compare_arithmetic();
        bit comp = 1;
        comp &= arithmetic_exp_result.valid == txn_out.result.valid;
        for (int i=0; i<RISCV_V_NUM_BYTES_DATA; i++) begin
            if (arithmetic_exp_result.valid[i]) begin
                comp &= arithmetic_exp_result.data.Byte[i] == txn_out.result.data.Byte[i];
            end
        end
        if (~arithmetic_in_txn.is_reduct) begin
            comp &= compare_flags(arithmetic_in_txn.osize, arithmetic_exp_result.valid);
        end
        if (comp) begin
            pass();
        end else begin
            `uvm_error(get_name(), $sformatf("Compare mismatch, actual.valid: 0x%0h, actual.data: 0x%0h, actual.zf: 0x%0h, actual.of: 0x%0h, actual.cf: 0x%0h, exp.valid: 0x%0h, exp.data: 0x%0h, exp.zf: 0x%0h, exp.of: 0x%0h, exp.cf: 0x%0h", txn_out.result.valid, txn_out.result.data, txn_out.zf, txn_out.of, txn_out.cf, arithmetic_exp_result.valid, arithmetic_exp_result.data, zf_exp, of_exp, cf_exp))
            fail();
        end
    endfunction: compare_arithmetic

    virtual function void compare_mask();
        riscv_v_mask_alu_out_seq_item mask_txn_out;
        bit comp = 1;

        if (!$cast(mask_txn_out, txn_out)) begin
            `uvm_fatal(get_name(), "Can't cast txn_out to mask_txn_out")
        end

        for (int i=0; i < RISCV_V_NUM_ELEMENTS_REG; i++) begin
            comp &= mask_exp_result[i]  == mask_txn_out.result_mask[i];
        end

        if (comp) begin
            pass();
        end else begin
            `uvm_error(get_name(), $sformatf("Compare mismatch, actual.data: 0x%0h, exp.data: 0x%0h", mask_txn_out.result_mask, mask_exp_result))
            fail();
        end
    endfunction: compare_mask

    virtual function void compare_permutation();
        riscv_v_permutation_alu_out_seq_item permutation_txn_out;
        bit comp = 1;
        if (!$cast(permutation_txn_out, txn_out)) begin
            `uvm_fatal(get_name(), "Can't cast txn_out to permutation_txn_out")
        end

        comp &= (permutation_exp_int_result       == permutation_txn_out.integer_data_out);
        comp &= (permutation_exp_vec_result.data  == permutation_txn_out.vector_data_out.data);
        comp &= (permutation_exp_vec_result.valid == permutation_txn_out.vector_data_out.valid);

        if (comp) begin
            pass();
        end else begin
            `uvm_error(get_name(), $sformatf("Compare mismatch, actual_int.data: 0x%0h, actual_vec.data: 0x%0h, actual_vec.valid: 0x%0h, exp_int.data: 0x%0h, exp_vec.data: 0x%0h, exp_vec.valid: 0x%0h", permutation_txn_out.integer_data_out, permutation_txn_out.vector_data_out.data, permutation_txn_out.vector_data_out.valid, permutation_exp_int_result, permutation_exp_vec_result.data, permutation_exp_vec_result.valid))
            fail();
        end

    endfunction: compare_permutation

    virtual function bit compare_flags(riscv_v_osize_e osize, riscv_v_valid_data_t valid);
        bit comp = 1;
        case (osize)
            OSIZE_8: begin
                for (int i=0; i<RISCV_V_NUM_BYTES_DATA; i++) begin
                    if (valid[i]) begin
                        comp &= zf_exp[i] == txn_out.zf[i];
                        comp &= cf_exp[i] == txn_out.cf[i];
                        comp &= of_exp[i] == txn_out.of[i];
                    end
                end
            end
            OSIZE_16: begin
                for (int i=0; i<RISCV_V_NUM_WORDS_DATA; i++) begin
                    if (valid[(i*2)+1]) begin
                        comp &= zf_exp[(i*2)+1] == txn_out.zf[(i*2)+1];
                        comp &= cf_exp[(i*2)+1] == txn_out.cf[(i*2)+1];
                        comp &= of_exp[(i*2)+1] == txn_out.of[(i*2)+1];
                    end
                end
            end
            OSIZE_32: begin
                for (int i=0; i<RISCV_V_NUM_DWORDS_DATA; i++) begin
                    if (valid[(i*4)+3]) begin
                        comp &= zf_exp[(i*4)+3] == txn_out.zf[(i*4)+3];
                        comp &= cf_exp[(i*4)+3] == txn_out.cf[(i*4)+3];
                        comp &= of_exp[(i*4)+3] == txn_out.of[(i*4)+3];
                    end
                end
            end
            OSIZE_64: begin
                for (int i=0; i<RISCV_V_NUM_QWORDS_DATA; i++) begin
                    if (valid[(i*8)+7]) begin
                        comp &= zf_exp[(i*8)+7] == txn_out.zf[(i*8)+7];
                        comp &= cf_exp[(i*8)+7] == txn_out.cf[(i*8)+7];
                        comp &= of_exp[(i*8)+7] == txn_out.of[(i*8)+7];
                    end
                end
            end
            OSIZE_128: begin
                for (int i=0; i<RISCV_V_NUM_DQWORDS_DATA; i++) begin
                    if (valid[(i*16)+15]) begin
                        comp &= zf_exp[(i*16)+15] == txn_out.zf[(i*16)+15];
                        comp &= cf_exp[(i*16)+15] == txn_out.cf[(i*16)+15];
                        comp &= of_exp[(i*16)+15] == txn_out.of[(i*16)+15];
                    end
                end
            end
            default: `uvm_fatal(get_name(), "Invalid osize in compare_flags()")
        endcase
        return comp;
    endfunction: compare_flags

    virtual function void calc_valid();
        logic_exp_result.valid = txn_in.srca.valid;
        arithmetic_exp_result.valid = txn_in.srca.valid;
    endfunction: calc_valid

    `include "riscv_v_alu_scbd_logic_ops.sv"
    `include "riscv_v_alu_scbd_arithmetic_ops.sv"
    `include "riscv_v_alu_scbd_mask_ops.sv"
    `include "riscv_v_alu_scbd_permutation_ops.sv"

endclass: riscv_v_alu_scbd

`endif // __RISCV_V_ALU_SCBD_SV__