module riscv_v_memory (
	clk,
	rst
);
	input wire clk;
	input wire rst;
endmodule
