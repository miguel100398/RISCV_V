//File: riscv_v_cpu_vredsum_test
//Author: Miguel Bucio
//Date: 10/02/24
//Description: RISC-V Vector CPU Reduction ADD Test

`ifndef __RISCV_V_CPU_VREDSUM_TEST_SV__
`define __RISCV_V_CPU_VREDSUM_TEST_SV__

class riscv_v_cpu_vredsum_test extends riscv_v_cpu_base_test;

    `uvm_component_utils(riscv_v_cpu_vredsum_test)

    function new(string name = "riscv_v_cpu_vredsum_test",uvm_component parent=null);
        super.new(name,parent);
        //Set Global variables
        NUM_TXN_BLOCK  = 50;
        SUPPORTS_MASK  = 1;
        NUM_OSIZES     = RISCV_V_NUM_VALID_OSIZES-1;
        NUM_FORMATS    = 1;
        TOTAL_BLOCKS   = NUM_FORMATS*NUM_OSIZES*(SUPPORTS_MASK+1);
        USE_RAND_START = 1'b0;
        USE_RAND_LEN   = 1'b1;
    endfunction : new

    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase);
    endfunction : build_phase

    virtual function void specific_bfm_cfg();
        //Instruction Fetch
        if_cfg.use_specific_instr   = 1'b1;
        if_cfg.use_specific_mode    = 1'b1;
        if_cfg.use_specific_vm      = 1'b1;
        if_cfg.specific_instr       = ADD_REDUCT;
        if_cfg.specific_mode        = OPIVV;
        if_cfg.specific_vm          = 1'b1;
        //Set Valid osizes for test
        valid_osizes = new[NUM_OSIZES];
        valid_osizes = '{OSIZE_8, OSIZE_16, OSIZE_32, OSIZE_64};
        //Set Valid formats for test
        valid_formats = new[NUM_FORMATS];
        valid_formats = '{OPMVV};
        //Dont update vstart
        cfg_wr_vstart = 1'b0;

    endfunction: specific_bfm_cfg

endclass: riscv_v_cpu_vredsum_test 

`endif //__RISCV_V_CPU_VREDSUM_TEST_SV__ 