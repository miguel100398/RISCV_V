//File: riscv_v_memory.sv
//Author: Miguel Bucio
//Date: 15/01/24
//Description: RISC-V Vector extension Memory Stage

module riscv_v_memory
import riscv_pkg::*, riscv_v_pkg::*;
(
    //Clocks and resets
    input  logic clk,
    input  logic rst
);

endmodule: riscv_v_memory