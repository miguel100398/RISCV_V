//File: riscv_v_alu_test_pkg.sv
//Author: Miguel Bucio
//Date: 11/02/24
//Description: RISC-V Vector ALU test package

package riscv_v_alu_test_pkg;
    import uvm_pkg::*; 
    import riscv_pkg::*;
    import riscv_v_pkg::*;
    import riscv_v_alu_agt_pkg::*;

    `include "uvm_macros.svh"
    import riscv_v_base_test_pkg::*;
    import riscv_v_base_alu_test_pkg::*;
    import riscv_v_arithmetic_alu_test_pkg::*;
    import riscv_v_logic_alu_test_pkg::*;
    import riscv_v_mask_alu_test_pkg::*;
    import riscv_v_permutation_alu_test_pkg::*;

endpackage: riscv_v_alu_test_pkg
