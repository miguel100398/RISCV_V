//Description: GPIO package, defines common types and parameters used by GPIO
//Author: Miguel Bucio miguel_angel_bucio@hotmail.com
//Date: 3/13/2022

package GPIO_pkg;

parameter GPIO_PORT_OUT_ADDR = 32'h10010024;
parameter GPIO_PORT_IN_ADDR  = 32'h10010028;

endpackage: GPIO_pkg