//File: riscv_v_test_pkg.sv
//Author: Miguel Bucio
//Date: 11/04/23
//Description: RISC-V Vector test package

package riscv_v_test_pkg;
    import riscv_v_pkg::*;
    import uvm_pkg::*;
    
    import riscv_v_alu_agt_pkg::*;

    
    `include "uvm_macros.svh"
    import riscv_v_base_test_pkg::*;
    import riscv_v_rf_test_pkg::*;
    import riscv_v_base_alu_test_pkg::*;
    import riscv_v_alu_test_pkg::*;
    import riscv_v_cpu_test_pkg::*;

endpackage: riscv_v_test_pkg