//File: riscv_v_base_test_pkg.sv
//Author: Miguel Bucio
//Date: 11/02/24
//Description: RISC-V Vector Base test package

package riscv_v_base_test_pkg;
    import uvm_pkg::*; 
    import riscv_pkg::*;
    import riscv_v_pkg::*;

    `include "uvm_macros.svh"
    `include "riscv_v_base_test.sv"

endpackage: riscv_v_base_test_pkg